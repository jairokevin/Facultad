LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all; 
USE IEEE.std_logic_unsigned.ALL; 

ENTITY signext IS
	GENERIC (N: INTEGER := 64);
	PORT (a: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			y: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0));               
END;
ARCHITECTURE synth of signext IS
BEGIN
	WITH a(31 DOWNTO 21) SELECT
		y <= STD_LOGIC_VECTOR(RESIZE(SIGNED(a(20 DOWNTO 12)), y'LENGTH)) 
				WHEN "11111000010" | "11111000000", --instruction type D
			 STD_LOGIC_VECTOR(RESIZE(SIGNED(a(23 DOWNTO 5)), y'LENGTH)) 
				WHEN "10110100000" | "10110100001" | "10110100010" | "10110100011" |
					  "10110100100" | "10110100101" | "10110100110" | "10110100111" | 
					  "10110101000" | "10110101001" | "10110101010" | "10110101011" |
					  "10110101100" | "10110101101" | "10110101110" | "10110101111" , --intruction type CB
			 STD_LOGIC_VECTOR(RESIZE(SIGNED(a(21 DOWNTO 10)), y'LENGTH))
				WHEN "10010001000" | "10010001001" , --instruction ADDI
			(OTHERS => '0') WHEN OTHERS;
				
END synth;	
